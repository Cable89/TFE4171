HDLC_packet test_message[10];

